
module ppi8255A(PortA,PortB,PortC,Re,Wr,Reset,A,Cs)




endmodule 